    assert false report "End of Testbench" severity FAILURE;
end process;
end block;
end architecture;